`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 12/04/2023 04:11:39 PM 
// Module Name: ALU
// Module Description :it takes 2 16 bit numbers and adds them 
//////////////////////////////////////////////////////////////////////////////////
module ALU (
input [15:0] A, P,
output reg [15:0] Result
);
assign Result = A + P; // addition

endmodule
