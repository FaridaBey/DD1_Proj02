`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/04/2023 04:11:39 PM
// Design Name: 
// Module Name: multiplier
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module multiplier(
    input  [7:0] multiplicand,
    input  [7:0] multiplier,
    input clk, reset,
    input load, enable, product_sel,
    output reg  [15:0] product,
    output  sign,
    output  zero_flag, b0 
);



endmodule
